----------------------------------------------------------------------------------
-- Company: Digilent Ro
-- Engineer: Tudor Armand Ciuleanu
-- 
-- Create Date:    10:51:31 02/28/2008 
-- Module Name:    LS1RefProj.vhd
-- Project Name: 	 LS1ReferenceProject
-- Tool versions:  Xilinx ISE 9.2
-- Description: This is the top module of the LS1 Reference Project. The 
--				SoundGenerator module and the Da2_controller module are instantiated
--				here.The sinus wave generated by the SoundGenerator module is sent to
--				the data1 input of the DA2_controller module. The SoundGenerator adds
--				together four sinus corresponding to different musical sounds(C, E, G, C)
--				A sound is added to the output if the coresponding bit returned by PmodLS1
--				HIGH.
--
-- Revision: 
-- Revision 0.01 - File Created
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity LS1RefProj is
    Port ( 	ck			: in STD_LOGIC;	--50 mhz clock input
			
			--LS1 signals	
				LSData 	: in  STD_LOGIC_VECTOR (3 downto 0); 
									
			--DA2 signals
				DAData 	: out  STD_LOGIC;				
				DAClk 	: out  STD_LOGIC;
				DASync 	: out  STD_LOGIC
				);
end LS1RefProj;

architecture Behavioral of LS1RefProj is

component DA2Component is
    Port ( 
	 --General usage
	   CLK      : in std_logic;	-- System Clock (50MHz)     
		RST		: in std_logic;
	 
	 --Pmod interface signals
      D1       : out std_logic;
	   D2		   : out std_logic;
		CLK_OUT	: out std_logic;
		nSYNC    : out std_logic;
		
	--User interface signals
	 	DATA1    : in std_logic_vector(11 downto 0);
		DATA2    : in std_logic_vector(11 downto 0);
	 	START	   : in std_logic; 
      DONE     : out std_logic 
		);
end component;

component SoundGenerator is
    Port ( ck 			: in  STD_LOGIC;
           LSData 	: in  STD_LOGIC_VECTOR (3 downto 0);
           SoundOut 	: out  STD_LOGIC_VECTOR (11 downto 0));
end component;

signal sync: STD_LOGIC;
signal sound: STD_LOGIC_VECTOR (11 downto 0);

begin

SoundGenerator_inst: SoundGenerator 
    Port Map( 
		ck 		=> ck	,
      LSData 	=> LSData,
      SoundOut => sound
		);	

DA2_inst: DA2Component
	port map (
		 --General usage
	   CLK 		=>  ck,
		RST		=>	 '0',
	 
	 --Pmod interface signals
      D1       =>	DAData,
	   D2		   =>	open,
		CLK_OUT	=> DAClk,
		nSYNC    => DASync,
		
	--User interface signals
	 	DATA1    =>	sound,	--sin wave from SoundGenerator
		DATA2    =>	"000000000000",
		--by connecting start and done together the da2
		--samples the data input at the highest rate possible 
	 	START	   => sync,		
      DONE     => sync
		);

end Behavioral;

